
// ハフマンテーブル
BitString y_dc_table[0:11];  // 輝度DCハフマンテーブル
BitString y_ac_table[0:255];  // 輝度ACハフマンテーブル
BitString cbcr_dc_table[0:11];  // 色差DCハフマンテーブル
BitString cbcr_ac_table[0:255];  // 色差ACハフマンテーブル

// ハフマンテーブル（Cコードに基づく全エントリ）
// 輝度DCハフマンテーブル（12エントリ）
//BitString y_dc_table[0:11];
initial begin
  y_dc_table[0]  = '{value: 16'h0006, length: 5'd3};
  y_dc_table[1]  = '{value: 16'h0005, length: 5'd3};
  y_dc_table[2]  = '{value: 16'h0003, length: 5'd3};
  y_dc_table[3]  = '{value: 16'h0002, length: 5'd3};
  y_dc_table[4]  = '{value: 16'h0000, length: 5'd3};
  y_dc_table[5]  = '{value: 16'h0001, length: 5'd3};
  y_dc_table[6]  = '{value: 16'h0004, length: 5'd3};
  y_dc_table[7]  = '{value: 16'h000e, length: 5'd4};
  y_dc_table[8]  = '{value: 16'h001e, length: 5'd5};
  y_dc_table[9]  = '{value: 16'h003e, length: 5'd6};
  y_dc_table[10] = '{value: 16'h007e, length: 5'd7};
  y_dc_table[11] = '{value: 16'h00fe, length: 5'd8};
end

// 輝度ACハフマンテーブル（162エントリ、CコードのStandard_AC_Luminance_Values）
//BitString y_ac_table[0:255];
initial begin
  y_ac_table[0]   = '{value: 16'h000a, length: 5'd4};
  y_ac_table[1]   = '{value: 16'h0000, length: 5'd2};
  y_ac_table[2]   = '{value: 16'h0001, length: 5'd2};
  y_ac_table[3]   = '{value: 16'h0004, length: 5'd3};
  y_ac_table[4]   = '{value: 16'h000b, length: 5'd4};
  y_ac_table[5]   = '{value: 16'h001a, length: 5'd5};
  y_ac_table[6]   = '{value: 16'h0078, length: 5'd7};
  y_ac_table[7]   = '{value: 16'h00f8, length: 5'd8};
  y_ac_table[8]   = '{value: 16'h03f6, length: 5'd10};
  y_ac_table[9]   = '{value: 16'hff82, length: 5'd16};
  y_ac_table[10]  = '{value: 16'hff83, length: 5'd16};
  y_ac_table[11]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[12]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[13]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[14]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[15]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[16]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[17]  = '{value: 16'h000c, length: 5'd4};
  y_ac_table[18]  = '{value: 16'h001b, length: 5'd5};
  y_ac_table[19]  = '{value: 16'h0079, length: 5'd7};
  y_ac_table[20]  = '{value: 16'h01f6, length: 5'd9};
  y_ac_table[21]  = '{value: 16'h07f6, length: 5'd11};
  y_ac_table[22]  = '{value: 16'hff84, length: 5'd16};
  y_ac_table[23]  = '{value: 16'hff85, length: 5'd16};
  y_ac_table[24]  = '{value: 16'hff86, length: 5'd16};
  y_ac_table[25]  = '{value: 16'hff87, length: 5'd16};
  y_ac_table[26]  = '{value: 16'hff88, length: 5'd16};
  y_ac_table[27]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[28]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[29]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[30]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[31]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[32]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[33]  = '{value: 16'h001c, length: 5'd5};
  y_ac_table[34]  = '{value: 16'h00f9, length: 5'd8};
  y_ac_table[35]  = '{value: 16'h03f7, length: 5'd10};
  y_ac_table[36]  = '{value: 16'h0ff4, length: 5'd12};
  y_ac_table[37]  = '{value: 16'hff89, length: 5'd16};
  y_ac_table[38]  = '{value: 16'hff8a, length: 5'd16};
  y_ac_table[39]  = '{value: 16'hff8b, length: 5'd16};
  y_ac_table[40]  = '{value: 16'hff8c, length: 5'd16};
  y_ac_table[41]  = '{value: 16'hff8d, length: 5'd16};
  y_ac_table[42]  = '{value: 16'hff8e, length: 5'd16};
  y_ac_table[43]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[44]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[45]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[46]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[47]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[48]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[49]  = '{value: 16'h003a, length: 5'd6};
  y_ac_table[50]  = '{value: 16'h01f7, length: 5'd9};
  y_ac_table[51]  = '{value: 16'h0ff5, length: 5'd12};
  y_ac_table[52]  = '{value: 16'hff8f, length: 5'd16};
  y_ac_table[53]  = '{value: 16'hff90, length: 5'd16};
  y_ac_table[54]  = '{value: 16'hff91, length: 5'd16};
  y_ac_table[55]  = '{value: 16'hff92, length: 5'd16};
  y_ac_table[56]  = '{value: 16'hff93, length: 5'd16};
  y_ac_table[57]  = '{value: 16'hff94, length: 5'd16};
  y_ac_table[58]  = '{value: 16'hff95, length: 5'd16};
  y_ac_table[59]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[60]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[61]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[62]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[63]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[64]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[65]  = '{value: 16'h003b, length: 5'd6};
  y_ac_table[66]  = '{value: 16'h03f8, length: 5'd10};
  y_ac_table[67]  = '{value: 16'hff96, length: 5'd16};
  y_ac_table[68]  = '{value: 16'hff97, length: 5'd16};
  y_ac_table[69]  = '{value: 16'hff98, length: 5'd16};
  y_ac_table[70]  = '{value: 16'hff99, length: 5'd16};
  y_ac_table[71]  = '{value: 16'hff9a, length: 5'd16};
  y_ac_table[72]  = '{value: 16'hff9b, length: 5'd16};
  y_ac_table[73]  = '{value: 16'hff9c, length: 5'd16};
  y_ac_table[74]  = '{value: 16'hff9d, length: 5'd16};
  y_ac_table[75]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[76]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[77]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[78]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[79]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[80]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[81]  = '{value: 16'h007a, length: 5'd7};
  y_ac_table[82]  = '{value: 16'h07f7, length: 5'd11};
  y_ac_table[83]  = '{value: 16'hff9e, length: 5'd16};
  y_ac_table[84]  = '{value: 16'hff9f, length: 5'd16};
  y_ac_table[85]  = '{value: 16'hffa0, length: 5'd16};
  y_ac_table[86]  = '{value: 16'hffa1, length: 5'd16};
  y_ac_table[87]  = '{value: 16'hffa2, length: 5'd16};
  y_ac_table[88]  = '{value: 16'hffa3, length: 5'd16};
  y_ac_table[89]  = '{value: 16'hffa4, length: 5'd16};
  y_ac_table[90]  = '{value: 16'hffa5, length: 5'd16};
  y_ac_table[91]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[92]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[93]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[94]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[95]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[96]  = '{value: 16'h0000, length: 5'd0};
  y_ac_table[97]  = '{value: 16'h007b, length: 5'd7};
  y_ac_table[98]  = '{value: 16'h0ff6, length: 5'd12};
  y_ac_table[99]  = '{value: 16'hffa6, length: 5'd16};
  y_ac_table[100] = '{value: 16'hffa7, length: 5'd16};
  y_ac_table[101] = '{value: 16'hffa8, length: 5'd16};
  y_ac_table[102] = '{value: 16'hffa9, length: 5'd16};
  y_ac_table[103] = '{value: 16'hffaa, length: 5'd16};
  y_ac_table[104] = '{value: 16'hffab, length: 5'd16};
  y_ac_table[105] = '{value: 16'hffac, length: 5'd16};
  y_ac_table[106] = '{value: 16'hffad, length: 5'd16};
  y_ac_table[107] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[108] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[109] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[110] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[111] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[112] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[113] = '{value: 16'h00fa, length: 5'd8};
  y_ac_table[114] = '{value: 16'h0ff7, length: 5'd12};
  y_ac_table[115] = '{value: 16'hffae, length: 5'd16};
  y_ac_table[116] = '{value: 16'hffaf, length: 5'd16};
  y_ac_table[117] = '{value: 16'hffb0, length: 5'd16};
  y_ac_table[118] = '{value: 16'hffb1, length: 5'd16};
  y_ac_table[119] = '{value: 16'hffb2, length: 5'd16};
  y_ac_table[120] = '{value: 16'hffb3, length: 5'd16};
  y_ac_table[121] = '{value: 16'hffb4, length: 5'd16};
  y_ac_table[122] = '{value: 16'hffb5, length: 5'd16};
  y_ac_table[123] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[124] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[125] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[126] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[127] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[128] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[129] = '{value: 16'h01f8, length: 5'd9};
  y_ac_table[130] = '{value: 16'h7fc0, length: 5'd15};
  y_ac_table[131] = '{value: 16'hffb6, length: 5'd16};
  y_ac_table[132] = '{value: 16'hffb7, length: 5'd16};
  y_ac_table[133] = '{value: 16'hffb8, length: 5'd16};
  y_ac_table[134] = '{value: 16'hffb9, length: 5'd16};
  y_ac_table[135] = '{value: 16'hffba, length: 5'd16};
  y_ac_table[136] = '{value: 16'hffbb, length: 5'd16};
  y_ac_table[137] = '{value: 16'hffbc, length: 5'd16};
  y_ac_table[138] = '{value: 16'hffbd, length: 5'd16};
  y_ac_table[139] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[140] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[141] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[142] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[143] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[144] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[145] = '{value: 16'h01f9, length: 5'd9};
  y_ac_table[146] = '{value: 16'hffbe, length: 5'd16};
  y_ac_table[147] = '{value: 16'hffbf, length: 5'd16};
  y_ac_table[148] = '{value: 16'hffc0, length: 5'd16};
  y_ac_table[149] = '{value: 16'hffc1, length: 5'd16};
  y_ac_table[150] = '{value: 16'hffc2, length: 5'd16};
  y_ac_table[151] = '{value: 16'hffc3, length: 5'd16};
  y_ac_table[152] = '{value: 16'hffc4, length: 5'd16};
  y_ac_table[153] = '{value: 16'hffc5, length: 5'd16};
  y_ac_table[154] = '{value: 16'hffc6, length: 5'd16};
  y_ac_table[155] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[156] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[157] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[158] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[159] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[160] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[161] = '{value: 16'h01fa, length: 5'd9};
  y_ac_table[162] = '{value: 16'hffc7, length: 5'd16};
  y_ac_table[163] = '{value: 16'hffc8, length: 5'd16};
  y_ac_table[164] = '{value: 16'hffc9, length: 5'd16};
  y_ac_table[165] = '{value: 16'hffca, length: 5'd16};
  y_ac_table[166] = '{value: 16'hffcb, length: 5'd16};
  y_ac_table[167] = '{value: 16'hffcc, length: 5'd16};
  y_ac_table[168] = '{value: 16'hffcd, length: 5'd16};
  y_ac_table[169] = '{value: 16'hffce, length: 5'd16};
  y_ac_table[170] = '{value: 16'hffcf, length: 5'd16};
  y_ac_table[171] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[172] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[173] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[174] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[175] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[176] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[177] = '{value: 16'h03f9, length: 5'd10};
  y_ac_table[178] = '{value: 16'hffd0, length: 5'd16};
  y_ac_table[179] = '{value: 16'hffd1, length: 5'd16};
  y_ac_table[180] = '{value: 16'hffd2, length: 5'd16};
  y_ac_table[181] = '{value: 16'hffd3, length: 5'd16};
  y_ac_table[182] = '{value: 16'hffd4, length: 5'd16};
  y_ac_table[183] = '{value: 16'hffd5, length: 5'd16};
  y_ac_table[184] = '{value: 16'hffd6, length: 5'd16};
  y_ac_table[185] = '{value: 16'hffd7, length: 5'd16};
  y_ac_table[186] = '{value: 16'hffd8, length: 5'd16};
  y_ac_table[187] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[188] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[189] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[190] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[191] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[192] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[193] = '{value: 16'h03fa, length: 5'd10};
  y_ac_table[194] = '{value: 16'hffd9, length: 5'd16};
  y_ac_table[195] = '{value: 16'hffda, length: 5'd16};
  y_ac_table[196] = '{value: 16'hffdb, length: 5'd16};
  y_ac_table[197] = '{value: 16'hffdc, length: 5'd16};
  y_ac_table[198] = '{value: 16'hffdd, length: 5'd16};
  y_ac_table[199] = '{value: 16'hffde, length: 5'd16};
  y_ac_table[200] = '{value: 16'hffdf, length: 5'd16};
  y_ac_table[201] = '{value: 16'hffe0, length: 5'd16};
  y_ac_table[202] = '{value: 16'hffe1, length: 5'd16};
  y_ac_table[203] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[204] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[205] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[206] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[207] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[208] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[209] = '{value: 16'h07f8, length: 5'd11};
  y_ac_table[210] = '{value: 16'hffe2, length: 5'd16};
  y_ac_table[211] = '{value: 16'hffe3, length: 5'd16};
  y_ac_table[212] = '{value: 16'hffe4, length: 5'd16};
  y_ac_table[213] = '{value: 16'hffe5, length: 5'd16};
  y_ac_table[214] = '{value: 16'hffe6, length: 5'd16};
  y_ac_table[215] = '{value: 16'hffe7, length: 5'd16};
  y_ac_table[216] = '{value: 16'hffe8, length: 5'd16};
  y_ac_table[217] = '{value: 16'hffe9, length: 5'd16};
  y_ac_table[218] = '{value: 16'hffea, length: 5'd16};
  y_ac_table[219] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[220] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[221] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[222] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[223] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[224] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[225] = '{value: 16'hffeb, length: 5'd16};
  y_ac_table[226] = '{value: 16'hffec, length: 5'd16};
  y_ac_table[227] = '{value: 16'hffed, length: 5'd16};
  y_ac_table[228] = '{value: 16'hffee, length: 5'd16};
  y_ac_table[229] = '{value: 16'hffef, length: 5'd16};
  y_ac_table[230] = '{value: 16'hfff0, length: 5'd16};
  y_ac_table[231] = '{value: 16'hfff1, length: 5'd16};
  y_ac_table[232] = '{value: 16'hfff2, length: 5'd16};
  y_ac_table[233] = '{value: 16'hfff3, length: 5'd16};
  y_ac_table[234] = '{value: 16'hfff4, length: 5'd16};
  y_ac_table[235] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[236] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[237] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[238] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[239] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[240] = '{value: 16'h07f9, length: 5'd11};
  y_ac_table[241] = '{value: 16'hfff5, length: 5'd16};
  y_ac_table[242] = '{value: 16'hfff6, length: 5'd16};
  y_ac_table[243] = '{value: 16'hfff7, length: 5'd16};
  y_ac_table[244] = '{value: 16'hfff8, length: 5'd16};
  y_ac_table[245] = '{value: 16'hfff9, length: 5'd16};
  y_ac_table[246] = '{value: 16'hfffa, length: 5'd16};
  y_ac_table[247] = '{value: 16'hfffb, length: 5'd16};
  y_ac_table[248] = '{value: 16'hfffc, length: 5'd16};
  y_ac_table[249] = '{value: 16'hfffd, length: 5'd16};
  y_ac_table[250] = '{value: 16'hfffe, length: 5'd16};
  y_ac_table[251] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[252] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[253] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[254] = '{value: 16'h0000, length: 5'd0};
  y_ac_table[255] = '{value: 16'h0000, length: 5'd0};
end

// 色差DCハフマンテーブル（12エントリ）
//BitString cbcr_dc_table[0:11];
initial begin
  cbcr_dc_table[0]  = '{value: 16'h0000, length: 5'd2};
  cbcr_dc_table[1]  = '{value: 16'h0001, length: 5'd2};
  cbcr_dc_table[2]  = '{value: 16'h0002, length: 5'd2};
  cbcr_dc_table[3]  = '{value: 16'h0006, length: 5'd3};
  cbcr_dc_table[4]  = '{value: 16'h000e, length: 5'd4};
  cbcr_dc_table[5]  = '{value: 16'h001e, length: 5'd5};
  cbcr_dc_table[6]  = '{value: 16'h003e, length: 5'd6};
  cbcr_dc_table[7]  = '{value: 16'h007e, length: 5'd7};
  cbcr_dc_table[8]  = '{value: 16'h00fe, length: 5'd8};
  cbcr_dc_table[9]  = '{value: 16'h01fe, length: 5'd9};
  cbcr_dc_table[10] = '{value: 16'h03fe, length: 5'd10};
  cbcr_dc_table[11] = '{value: 16'h07fe, length: 5'd11};
end

// 色差ACハフマンテーブル（162エントリ、CコードのStandard_AC_Chrominance_Values）
//BitString cbcr_ac_table[0:255];
initial begin
  cbcr_ac_table[0]   = '{value: 16'h0000, length: 5'd2};
  cbcr_ac_table[1]   = '{value: 16'h0001, length: 5'd2};
  cbcr_ac_table[2]   = '{value: 16'h0004, length: 5'd3};
  cbcr_ac_table[3]   = '{value: 16'h000a, length: 5'd4};
  cbcr_ac_table[4]   = '{value: 16'h0018, length: 5'd5};
  cbcr_ac_table[5]   = '{value: 16'h0019, length: 5'd5};
  cbcr_ac_table[6]   = '{value: 16'h0038, length: 5'd6};
  cbcr_ac_table[7]   = '{value: 16'h0078, length: 5'd7};
  cbcr_ac_table[8]   = '{value: 16'h01f4, length: 5'd9};
  cbcr_ac_table[9]   = '{value: 16'h03f6, length: 5'd10};
  cbcr_ac_table[10]  = '{value: 16'h0ff4, length: 5'd12};
  cbcr_ac_table[11]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[12]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[13]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[14]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[15]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[16]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[17]  = '{value: 16'h000b, length: 5'd4};
  cbcr_ac_table[18]  = '{value: 16'h0039, length: 5'd6};
  cbcr_ac_table[19]  = '{value: 16'h00f6, length: 5'd8};
  cbcr_ac_table[20]  = '{value: 16'h01f5, length: 5'd9};
  cbcr_ac_table[21]  = '{value: 16'h07f6, length: 5'd11};
  cbcr_ac_table[22]  = '{value: 16'h0ff5, length: 5'd12};
  cbcr_ac_table[23]  = '{value: 16'hff88, length: 5'd16};
  cbcr_ac_table[24]  = '{value: 16'hff89, length: 5'd16};
  cbcr_ac_table[25]  = '{value: 16'hff8a, length: 5'd16};
  cbcr_ac_table[26]  = '{value: 16'hff8b, length: 5'd16};
  cbcr_ac_table[27]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[28]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[29]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[30]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[31]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[32]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[33]  = '{value: 16'h001a, length: 5'd5};
  cbcr_ac_table[34]  = '{value: 16'h00f7, length: 5'd8};
  cbcr_ac_table[35]  = '{value: 16'h03f7, length: 5'd10};
  cbcr_ac_table[36]  = '{value: 16'h0ff6, length: 5'd12};
  cbcr_ac_table[37]  = '{value: 16'h7fc2, length: 5'd15};
  cbcr_ac_table[38]  = '{value: 16'hff8c, length: 5'd16};
  cbcr_ac_table[39]  = '{value: 16'hff8d, length: 5'd16};
  cbcr_ac_table[40]  = '{value: 16'hff8e, length: 5'd16};
  cbcr_ac_table[41]  = '{value: 16'hff8f, length: 5'd16};
  cbcr_ac_table[42]  = '{value: 16'hff90, length: 5'd16};
  cbcr_ac_table[43]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[44]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[45]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[46]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[47]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[48]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[49]  = '{value: 16'h001b, length: 5'd5};
  cbcr_ac_table[50]  = '{value: 16'h00f8, length: 5'd8};
  cbcr_ac_table[51]  = '{value: 16'h03f8, length: 5'd10};
  cbcr_ac_table[52]  = '{value: 16'h0ff7, length: 5'd12};
  cbcr_ac_table[53]  = '{value: 16'hff91, length: 5'd16};
  cbcr_ac_table[54]  = '{value: 16'hff92, length: 5'd16};
  cbcr_ac_table[55]  = '{value: 16'hff93, length: 5'd16};
  cbcr_ac_table[56]  = '{value: 16'hff94, length: 5'd16};
  cbcr_ac_table[57]  = '{value: 16'hff95, length: 5'd16};
  cbcr_ac_table[58]  = '{value: 16'hff96, length: 5'd16};
  cbcr_ac_table[59]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[60]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[61]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[62]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[63]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[64]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[65]  = '{value: 16'h003a, length: 5'd6};
  cbcr_ac_table[66]  = '{value: 16'h01f6, length: 5'd9};
  cbcr_ac_table[67]  = '{value: 16'hff97, length: 5'd16};
  cbcr_ac_table[68]  = '{value: 16'hff98, length: 5'd16};
  cbcr_ac_table[69]  = '{value: 16'hff99, length: 5'd16};
  cbcr_ac_table[70]  = '{value: 16'hff9a, length: 5'd16};
  cbcr_ac_table[71]  = '{value: 16'hff9b, length: 5'd16};
  cbcr_ac_table[72]  = '{value: 16'hff9c, length: 5'd16};
  cbcr_ac_table[73]  = '{value: 16'hff9d, length: 5'd16};
  cbcr_ac_table[74]  = '{value: 16'hff9e, length: 5'd16};
  cbcr_ac_table[75]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[76]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[77]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[78]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[79]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[80]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[81]  = '{value: 16'h003b, length: 5'd6};
  cbcr_ac_table[82]  = '{value: 16'h03f9, length: 5'd10};
  cbcr_ac_table[83]  = '{value: 16'hff9f, length: 5'd16};
  cbcr_ac_table[84]  = '{value: 16'hffa0, length: 5'd16};
  cbcr_ac_table[85]  = '{value: 16'hffa1, length: 5'd16};
  cbcr_ac_table[86]  = '{value: 16'hffa2, length: 5'd16};
  cbcr_ac_table[87]  = '{value: 16'hffa3, length: 5'd16};
  cbcr_ac_table[88]  = '{value: 16'hffa4, length: 5'd16};
  cbcr_ac_table[89]  = '{value: 16'hffa5, length: 5'd16};
  cbcr_ac_table[90]  = '{value: 16'hffa6, length: 5'd16};
  cbcr_ac_table[91]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[92]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[93]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[94]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[95]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[96]  = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[97]  = '{value: 16'h0079, length: 5'd7};
  cbcr_ac_table[98]  = '{value: 16'h07f7, length: 5'd11};
  cbcr_ac_table[99]  = '{value: 16'hffa7, length: 5'd16};
  cbcr_ac_table[100] = '{value: 16'hffa8, length: 5'd16};
  cbcr_ac_table[101] = '{value: 16'hffa9, length: 5'd16};
  cbcr_ac_table[102] = '{value: 16'hffaa, length: 5'd16};
  cbcr_ac_table[103] = '{value: 16'hffab, length: 5'd16};
  cbcr_ac_table[104] = '{value: 16'hffac, length: 5'd16};
  cbcr_ac_table[105] = '{value: 16'hffad, length: 5'd16};
  cbcr_ac_table[106] = '{value: 16'hffae, length: 5'd16};
  cbcr_ac_table[107] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[108] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[109] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[110] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[111] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[112] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[113] = '{value: 16'h007a, length: 5'd7};
  cbcr_ac_table[114] = '{value: 16'h07f8, length: 5'd11};
  cbcr_ac_table[115] = '{value: 16'hffaf, length: 5'd16};
  cbcr_ac_table[116] = '{value: 16'hffb0, length: 5'd16};
  cbcr_ac_table[117] = '{value: 16'hffb1, length: 5'd16};
  cbcr_ac_table[118] = '{value: 16'hffb2, length: 5'd16};
  cbcr_ac_table[119] = '{value: 16'hffb3, length: 5'd16};
  cbcr_ac_table[120] = '{value: 16'hffb4, length: 5'd16};
  cbcr_ac_table[121] = '{value: 16'hffb5, length: 5'd16};
  cbcr_ac_table[122] = '{value: 16'hffb6, length: 5'd16};
  cbcr_ac_table[123] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[124] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[125] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[126] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[127] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[128] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[129] = '{value: 16'h00f9, length: 5'd8};
  cbcr_ac_table[130] = '{value: 16'hffb7, length: 5'd16};
  cbcr_ac_table[131] = '{value: 16'hffb8, length: 5'd16};
  cbcr_ac_table[132] = '{value: 16'hffb9, length: 5'd16};
  cbcr_ac_table[133] = '{value: 16'hffba, length: 5'd16};
  cbcr_ac_table[134] = '{value: 16'hffbb, length: 5'd16};
  cbcr_ac_table[135] = '{value: 16'hffbc, length: 5'd16};
  cbcr_ac_table[136] = '{value: 16'hffbd, length: 5'd16};
  cbcr_ac_table[137] = '{value: 16'hffbe, length: 5'd16};
  cbcr_ac_table[138] = '{value: 16'hffbf, length: 5'd16};
  cbcr_ac_table[139] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[140] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[141] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[142] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[143] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[144] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[145] = '{value: 16'h01f7, length: 5'd9};
  cbcr_ac_table[146] = '{value: 16'hffc0, length: 5'd16};
  cbcr_ac_table[147] = '{value: 16'hffc1, length: 5'd16};
  cbcr_ac_table[148] = '{value: 16'hffc2, length: 5'd16};
  cbcr_ac_table[149] = '{value: 16'hffc3, length: 5'd16};
  cbcr_ac_table[150] = '{value: 16'hffc4, length: 5'd16};
  cbcr_ac_table[151] = '{value: 16'hffc5, length: 5'd16};
  cbcr_ac_table[152] = '{value: 16'hffc6, length: 5'd16};
  cbcr_ac_table[153] = '{value: 16'hffc7, length: 5'd16};
  cbcr_ac_table[154] = '{value: 16'hffc8, length: 5'd16};
  cbcr_ac_table[155] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[156] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[157] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[158] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[159] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[160] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[161] = '{value: 16'h01f8, length: 5'd9};
  cbcr_ac_table[162] = '{value: 16'hffc9, length: 5'd16};
  cbcr_ac_table[163] = '{value: 16'hffca, length: 5'd16};
  cbcr_ac_table[164] = '{value: 16'hffcb, length: 5'd16};
  cbcr_ac_table[165] = '{value: 16'hffcc, length: 5'd16};
  cbcr_ac_table[166] = '{value: 16'hffcd, length: 5'd16};
  cbcr_ac_table[167] = '{value: 16'hffce, length: 5'd16};
  cbcr_ac_table[168] = '{value: 16'hffcf, length: 5'd16};
  cbcr_ac_table[169] = '{value: 16'hffd0, length: 5'd16};
  cbcr_ac_table[170] = '{value: 16'hffd1, length: 5'd16};
  cbcr_ac_table[171] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[172] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[173] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[174] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[175] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[176] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[177] = '{value: 16'h01f9, length: 5'd9};
  cbcr_ac_table[178] = '{value: 16'hffd2, length: 5'd16};
  cbcr_ac_table[179] = '{value: 16'hffd3, length: 5'd16};
  cbcr_ac_table[180] = '{value: 16'hffd4, length: 5'd16};
  cbcr_ac_table[181] = '{value: 16'hffd5, length: 5'd16};
  cbcr_ac_table[182] = '{value: 16'hffd6, length: 5'd16};
  cbcr_ac_table[183] = '{value: 16'hffd7, length: 5'd16};
  cbcr_ac_table[184] = '{value: 16'hffd8, length: 5'd16};
  cbcr_ac_table[185] = '{value: 16'hffd9, length: 5'd16};
  cbcr_ac_table[186] = '{value: 16'hffda, length: 5'd16};
  cbcr_ac_table[187] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[188] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[189] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[190] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[191] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[192] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[193] = '{value: 16'h01fa, length: 5'd9};
  cbcr_ac_table[194] = '{value: 16'hffdb, length: 5'd16};
  cbcr_ac_table[195] = '{value: 16'hffdc, length: 5'd16};
  cbcr_ac_table[196] = '{value: 16'hffdd, length: 5'd16};
  cbcr_ac_table[197] = '{value: 16'hffde, length: 5'd16};
  cbcr_ac_table[198] = '{value: 16'hffdf, length: 5'd16};
  cbcr_ac_table[199] = '{value: 16'hffe0, length: 5'd16};
  cbcr_ac_table[200] = '{value: 16'hffe1, length: 5'd16};
  cbcr_ac_table[201] = '{value: 16'hffe2, length: 5'd16};
  cbcr_ac_table[202] = '{value: 16'hffe3, length: 5'd16};
  cbcr_ac_table[203] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[204] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[205] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[206] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[207] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[208] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[209] = '{value: 16'h07f9, length: 5'd11};
  cbcr_ac_table[210] = '{value: 16'hffe4, length: 5'd16};
  cbcr_ac_table[211] = '{value: 16'hffe5, length: 5'd16};
  cbcr_ac_table[212] = '{value: 16'hffe6, length: 5'd16};
  cbcr_ac_table[213] = '{value: 16'hffe7, length: 5'd16};
  cbcr_ac_table[214] = '{value: 16'hffe8, length: 5'd16};
  cbcr_ac_table[215] = '{value: 16'hffe9, length: 5'd16};
  cbcr_ac_table[216] = '{value: 16'hffea, length: 5'd16};
  cbcr_ac_table[217] = '{value: 16'hffeb, length: 5'd16};
  cbcr_ac_table[218] = '{value: 16'hffec, length: 5'd16};
  cbcr_ac_table[219] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[220] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[221] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[222] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[223] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[224] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[225] = '{value: 16'h3fe0, length: 5'd14};
  cbcr_ac_table[226] = '{value: 16'hffed, length: 5'd16};
  cbcr_ac_table[227] = '{value: 16'hffee, length: 5'd16};
  cbcr_ac_table[228] = '{value: 16'hffef, length: 5'd16};
  cbcr_ac_table[229] = '{value: 16'hfff0, length: 5'd16};
  cbcr_ac_table[230] = '{value: 16'hfff1, length: 5'd16};
  cbcr_ac_table[231] = '{value: 16'hfff2, length: 5'd16};
  cbcr_ac_table[232] = '{value: 16'hfff3, length: 5'd16};
  cbcr_ac_table[233] = '{value: 16'hfff4, length: 5'd16};
  cbcr_ac_table[234] = '{value: 16'hfff5, length: 5'd16};
  cbcr_ac_table[235] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[236] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[237] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[238] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[239] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[240] = '{value: 16'h03fa, length: 5'd10};
  cbcr_ac_table[241] = '{value: 16'h7fc3, length: 5'd15};
  cbcr_ac_table[242] = '{value: 16'hfff6, length: 5'd16};
  cbcr_ac_table[243] = '{value: 16'hfff7, length: 5'd16};
  cbcr_ac_table[244] = '{value: 16'hfff8, length: 5'd16};
  cbcr_ac_table[245] = '{value: 16'hfff9, length: 5'd16};
  cbcr_ac_table[246] = '{value: 16'hfffa, length: 5'd16};
  cbcr_ac_table[247] = '{value: 16'hfffb, length: 5'd16};
  cbcr_ac_table[248] = '{value: 16'hfffc, length: 5'd16};
  cbcr_ac_table[249] = '{value: 16'hfffd, length: 5'd16};
  cbcr_ac_table[250] = '{value: 16'hfffe, length: 5'd16};
  cbcr_ac_table[251] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[252] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[253] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[254] = '{value: 16'h0000, length: 5'd0};
  cbcr_ac_table[255] = '{value: 16'h0000, length: 5'd0};
end
