
localparam signed [7:0] LUMA_QUANT_TABLE[0:63] = '{
    12,
    8,
    9,
    11,
    9,
    8,
    12,
    11,
    10,
    11,
    14,
    13,
    12,
    14,
    18,
    30,
    20,
    18,
    17,
    17,
    18,
    37,
    26,
    28,
    22,
    30,
    44,
    38,
    46,
    45,
    43,
    38,
    42,
    41,
    48,
    54,
    69,
    59,
    48,
    51,
    65,
    52,
    41,
    42,
    60,
    82,
    61,
    65,
    71,
    74,
    77,
    78,
    77,
    47,
    58,
    85,
    91,
    84,
    75,
    90,
    69,
    76,
    77,
    74
};

localparam signed [7:0] CHROMA_QUANT_TABLE[0:63] = '{
    13,
    14,
    14,
    18,
    16,
    18,
    35,
    20,
    20,
    35,
    74,
    50,
    42,
    50,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74,
    74
};
