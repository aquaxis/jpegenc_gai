// コサインテーブル（変更なし）
localparam logic signed [15:0] COS_TABLE[8][8] = '{
    '{16384, 16069, 15137, 13573, 11585, 9102, 6270, 3196},
    '{16384, 13573, 6270, -3196, -11585, -16069, -15137, -9102},
    '{16384, 9102, -6270, -16069, -11585, 3196, 15137, 13573},
    '{16384, 3196, -15137, -9102, 11585, 13573, -6270, -16069},
    '{16384, -3196, -15137, 9102, 11585, -13573, -6270, 16069},
    '{16384, -9102, -6270, 16069, -11585, -3196, 15137, -13573},
    '{16384, -13573, 6270, 3196, -11585, 16069, -15137, 9102},
    '{16384, -16069, 15137, -13573, 11585, -9102, 6270, -3196}
};
