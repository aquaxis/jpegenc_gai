// JPEGヘッダ（CコードのJpegEncoder_write_jpeg_headerを参考）
`define HEADER_SIZE 607
logic [7:0] header[0:606];

initial begin
  header[0]   = 8'hFF;
  header[1]   = 8'hD8;
  header[2]   = 8'hFF;
  header[3]   = 8'hE0;
  header[4]   = 8'h00;
  header[5]   = 8'h10;
  header[6]   = 8'h4A;
  header[7]   = 8'h46;
  header[8]   = 8'h49;
  header[9]   = 8'h46;
  header[10]  = 8'h00;
  header[11]  = 8'h01;
  header[12]  = 8'h01;
  header[13]  = 8'h00;
  header[14]  = 8'h00;
  header[15]  = 8'h01;
  header[16]  = 8'h00;
  header[17]  = 8'h01;
  header[18]  = 8'h00;
  header[19]  = 8'h00;
  header[20]  = 8'hFF;
  header[21]  = 8'hDB;
  header[22]  = 8'h00;
  header[23]  = 8'h84;
  header[24]  = 8'h00;
  header[25]  = 8'h0C;
  header[26]  = 8'h08;
  header[27]  = 8'h09;
  header[28]  = 8'h0B;
  header[29]  = 8'h09;
  header[30]  = 8'h08;
  header[31]  = 8'h0C;
  header[32]  = 8'h0B;
  header[33]  = 8'h0A;
  header[34]  = 8'h0B;
  header[35]  = 8'h0E;
  header[36]  = 8'h0D;
  header[37]  = 8'h0C;
  header[38]  = 8'h0E;
  header[39]  = 8'h12;
  header[40]  = 8'h1E;
  header[41]  = 8'h14;
  header[42]  = 8'h12;
  header[43]  = 8'h11;
  header[44]  = 8'h11;
  header[45]  = 8'h12;
  header[46]  = 8'h25;
  header[47]  = 8'h1A;
  header[48]  = 8'h1C;
  header[49]  = 8'h16;
  header[50]  = 8'h1E;
  header[51]  = 8'h2C;
  header[52]  = 8'h26;
  header[53]  = 8'h2E;
  header[54]  = 8'h2D;
  header[55]  = 8'h2B;
  header[56]  = 8'h26;
  header[57]  = 8'h2A;
  header[58]  = 8'h29;
  header[59]  = 8'h30;
  header[60]  = 8'h36;
  header[61]  = 8'h45;
  header[62]  = 8'h3B;
  header[63]  = 8'h30;
  header[64]  = 8'h33;
  header[65]  = 8'h41;
  header[66]  = 8'h34;
  header[67]  = 8'h29;
  header[68]  = 8'h2A;
  header[69]  = 8'h3C;
  header[70]  = 8'h52;
  header[71]  = 8'h3D;
  header[72]  = 8'h41;
  header[73]  = 8'h47;
  header[74]  = 8'h4A;
  header[75]  = 8'h4D;
  header[76]  = 8'h4E;
  header[77]  = 8'h4D;
  header[78]  = 8'h2F;
  header[79]  = 8'h3A;
  header[80]  = 8'h55;
  header[81]  = 8'h5B;
  header[82]  = 8'h54;
  header[83]  = 8'h4B;
  header[84]  = 8'h5A;
  header[85]  = 8'h45;
  header[86]  = 8'h4C;
  header[87]  = 8'h4D;
  header[88]  = 8'h4A;
  header[89]  = 8'h01;
  header[90]  = 8'h0D;
  header[91]  = 8'h0E;
  header[92]  = 8'h0E;
  header[93]  = 8'h12;
  header[94]  = 8'h10;
  header[95]  = 8'h12;
  header[96]  = 8'h23;
  header[97]  = 8'h14;
  header[98]  = 8'h14;
  header[99]  = 8'h23;
  header[100] = 8'h4A;
  header[101] = 8'h32;
  header[102] = 8'h2A;
  header[103] = 8'h32;
  header[104] = 8'h4A;
  header[105] = 8'h4A;
  header[106] = 8'h4A;
  header[107] = 8'h4A;
  header[108] = 8'h4A;
  header[109] = 8'h4A;
  header[110] = 8'h4A;
  header[111] = 8'h4A;
  header[112] = 8'h4A;
  header[113] = 8'h4A;
  header[114] = 8'h4A;
  header[115] = 8'h4A;
  header[116] = 8'h4A;
  header[117] = 8'h4A;
  header[118] = 8'h4A;
  header[119] = 8'h4A;
  header[120] = 8'h4A;
  header[121] = 8'h4A;
  header[122] = 8'h4A;
  header[123] = 8'h4A;
  header[124] = 8'h4A;
  header[125] = 8'h4A;
  header[126] = 8'h4A;
  header[127] = 8'h4A;
  header[128] = 8'h4A;
  header[129] = 8'h4A;
  header[130] = 8'h4A;
  header[131] = 8'h4A;
  header[132] = 8'h4A;
  header[133] = 8'h4A;
  header[134] = 8'h4A;
  header[135] = 8'h4A;
  header[136] = 8'h4A;
  header[137] = 8'h4A;
  header[138] = 8'h4A;
  header[139] = 8'h4A;
  header[140] = 8'h4A;
  header[141] = 8'h4A;
  header[142] = 8'h4A;
  header[143] = 8'h4A;
  header[144] = 8'h4A;
  header[145] = 8'h4A;
  header[146] = 8'h4A;
  header[147] = 8'h4A;
  header[148] = 8'h4A;
  header[149] = 8'h4A;
  header[150] = 8'h4A;
  header[151] = 8'h4A;
  header[152] = 8'h4A;
  header[153] = 8'h4A;
  header[154] = 8'hFF;
  header[155] = 8'hC0;
  header[156] = 8'h00;
  header[157] = 8'h11;
  header[158] = 8'h08;
  header[159] = 8'h01;
  header[160] = 8'hE0;
  header[161] = 8'h02;
  header[162] = 8'h80;
  header[163] = 8'h03;
  header[164] = 8'h01;
  header[165] = 8'h22;
  header[166] = 8'h00;
  header[167] = 8'h02;
  header[168] = 8'h11;
  header[169] = 8'h01;
  header[170] = 8'h03;
  header[171] = 8'h11;
  header[172] = 8'h01;
  header[173] = 8'hFF;
  header[174] = 8'hC4;
  header[175] = 8'h01;
  header[176] = 8'hA2;
  header[177] = 8'h00;
  header[178] = 8'h00;
  header[179] = 8'h00;
  header[180] = 8'h07;
  header[181] = 8'h01;
  header[182] = 8'h01;
  header[183] = 8'h01;
  header[184] = 8'h01;
  header[185] = 8'h01;
  header[186] = 8'h00;
  header[187] = 8'h00;
  header[188] = 8'h00;
  header[189] = 8'h00;
  header[190] = 8'h00;
  header[191] = 8'h00;
  header[192] = 8'h00;
  header[193] = 8'h00;
  header[194] = 8'h04;
  header[195] = 8'h05;
  header[196] = 8'h03;
  header[197] = 8'h02;
  header[198] = 8'h06;
  header[199] = 8'h01;
  header[200] = 8'h00;
  header[201] = 8'h07;
  header[202] = 8'h08;
  header[203] = 8'h09;
  header[204] = 8'h0A;
  header[205] = 8'h0B;
  header[206] = 8'h10;
  header[207] = 8'h00;
  header[208] = 8'h02;
  header[209] = 8'h01;
  header[210] = 8'h03;
  header[211] = 8'h03;
  header[212] = 8'h02;
  header[213] = 8'h04;
  header[214] = 8'h03;
  header[215] = 8'h05;
  header[216] = 8'h05;
  header[217] = 8'h04;
  header[218] = 8'h04;
  header[219] = 8'h00;
  header[220] = 8'h00;
  header[221] = 8'h01;
  header[222] = 8'h7D;
  header[223] = 8'h01;
  header[224] = 8'h02;
  header[225] = 8'h03;
  header[226] = 8'h00;
  header[227] = 8'h04;
  header[228] = 8'h11;
  header[229] = 8'h05;
  header[230] = 8'h12;
  header[231] = 8'h21;
  header[232] = 8'h31;
  header[233] = 8'h41;
  header[234] = 8'h06;
  header[235] = 8'h13;
  header[236] = 8'h51;
  header[237] = 8'h61;
  header[238] = 8'h07;
  header[239] = 8'h22;
  header[240] = 8'h71;
  header[241] = 8'h14;
  header[242] = 8'h32;
  header[243] = 8'h81;
  header[244] = 8'h91;
  header[245] = 8'hA1;
  header[246] = 8'h08;
  header[247] = 8'h23;
  header[248] = 8'h42;
  header[249] = 8'hB1;
  header[250] = 8'hC1;
  header[251] = 8'h15;
  header[252] = 8'h52;
  header[253] = 8'hD1;
  header[254] = 8'hF0;
  header[255] = 8'h24;
  header[256] = 8'h33;
  header[257] = 8'h62;
  header[258] = 8'h72;
  header[259] = 8'h82;
  header[260] = 8'h09;
  header[261] = 8'h0A;
  header[262] = 8'h16;
  header[263] = 8'h17;
  header[264] = 8'h18;
  header[265] = 8'h19;
  header[266] = 8'h1A;
  header[267] = 8'h25;
  header[268] = 8'h26;
  header[269] = 8'h27;
  header[270] = 8'h28;
  header[271] = 8'h29;
  header[272] = 8'h2A;
  header[273] = 8'h34;
  header[274] = 8'h35;
  header[275] = 8'h36;
  header[276] = 8'h37;
  header[277] = 8'h38;
  header[278] = 8'h39;
  header[279] = 8'h3A;
  header[280] = 8'h43;
  header[281] = 8'h44;
  header[282] = 8'h45;
  header[283] = 8'h46;
  header[284] = 8'h47;
  header[285] = 8'h48;
  header[286] = 8'h49;
  header[287] = 8'h4A;
  header[288] = 8'h53;
  header[289] = 8'h54;
  header[290] = 8'h55;
  header[291] = 8'h56;
  header[292] = 8'h57;
  header[293] = 8'h58;
  header[294] = 8'h59;
  header[295] = 8'h5A;
  header[296] = 8'h63;
  header[297] = 8'h64;
  header[298] = 8'h65;
  header[299] = 8'h66;
  header[300] = 8'h67;
  header[301] = 8'h68;
  header[302] = 8'h69;
  header[303] = 8'h6A;
  header[304] = 8'h73;
  header[305] = 8'h74;
  header[306] = 8'h75;
  header[307] = 8'h76;
  header[308] = 8'h77;
  header[309] = 8'h78;
  header[310] = 8'h79;
  header[311] = 8'h7A;
  header[312] = 8'h83;
  header[313] = 8'h84;
  header[314] = 8'h85;
  header[315] = 8'h86;
  header[316] = 8'h87;
  header[317] = 8'h88;
  header[318] = 8'h89;
  header[319] = 8'h8A;
  header[320] = 8'h92;
  header[321] = 8'h93;
  header[322] = 8'h94;
  header[323] = 8'h95;
  header[324] = 8'h96;
  header[325] = 8'h97;
  header[326] = 8'h98;
  header[327] = 8'h99;
  header[328] = 8'h9A;
  header[329] = 8'hA2;
  header[330] = 8'hA3;
  header[331] = 8'hA4;
  header[332] = 8'hA5;
  header[333] = 8'hA6;
  header[334] = 8'hA7;
  header[335] = 8'hA8;
  header[336] = 8'hA9;
  header[337] = 8'hAA;
  header[338] = 8'hB2;
  header[339] = 8'hB3;
  header[340] = 8'hB4;
  header[341] = 8'hB5;
  header[342] = 8'hB6;
  header[343] = 8'hB7;
  header[344] = 8'hB8;
  header[345] = 8'hB9;
  header[346] = 8'hBA;
  header[347] = 8'hC2;
  header[348] = 8'hC3;
  header[349] = 8'hC4;
  header[350] = 8'hC5;
  header[351] = 8'hC6;
  header[352] = 8'hC7;
  header[353] = 8'hC8;
  header[354] = 8'hC9;
  header[355] = 8'hCA;
  header[356] = 8'hD2;
  header[357] = 8'hD3;
  header[358] = 8'hD4;
  header[359] = 8'hD5;
  header[360] = 8'hD6;
  header[361] = 8'hD7;
  header[362] = 8'hD8;
  header[363] = 8'hD9;
  header[364] = 8'hDA;
  header[365] = 8'hE1;
  header[366] = 8'hE2;
  header[367] = 8'hE3;
  header[368] = 8'hE4;
  header[369] = 8'hE5;
  header[370] = 8'hE6;
  header[371] = 8'hE7;
  header[372] = 8'hE8;
  header[373] = 8'hE9;
  header[374] = 8'hEA;
  header[375] = 8'hF1;
  header[376] = 8'hF2;
  header[377] = 8'hF3;
  header[378] = 8'hF4;
  header[379] = 8'hF5;
  header[380] = 8'hF6;
  header[381] = 8'hF7;
  header[382] = 8'hF8;
  header[383] = 8'hF9;
  header[384] = 8'hFA;
  header[385] = 8'h01;
  header[386] = 8'h00;
  header[387] = 8'h03;
  header[388] = 8'h01;
  header[389] = 8'h01;
  header[390] = 8'h01;
  header[391] = 8'h01;
  header[392] = 8'h01;
  header[393] = 8'h01;
  header[394] = 8'h01;
  header[395] = 8'h01;
  header[396] = 8'h01;
  header[397] = 8'h00;
  header[398] = 8'h00;
  header[399] = 8'h00;
  header[400] = 8'h00;
  header[401] = 8'h00;
  header[402] = 8'h00;
  header[403] = 8'h01;
  header[404] = 8'h02;
  header[405] = 8'h03;
  header[406] = 8'h04;
  header[407] = 8'h05;
  header[408] = 8'h06;
  header[409] = 8'h07;
  header[410] = 8'h08;
  header[411] = 8'h09;
  header[412] = 8'h0A;
  header[413] = 8'h0B;
  header[414] = 8'h11;
  header[415] = 8'h00;
  header[416] = 8'h02;
  header[417] = 8'h01;
  header[418] = 8'h02;
  header[419] = 8'h04;
  header[420] = 8'h04;
  header[421] = 8'h03;
  header[422] = 8'h04;
  header[423] = 8'h07;
  header[424] = 8'h05;
  header[425] = 8'h04;
  header[426] = 8'h04;
  header[427] = 8'h00;
  header[428] = 8'h01;
  header[429] = 8'h02;
  header[430] = 8'h77;
  header[431] = 8'h00;
  header[432] = 8'h01;
  header[433] = 8'h02;
  header[434] = 8'h03;
  header[435] = 8'h11;
  header[436] = 8'h04;
  header[437] = 8'h05;
  header[438] = 8'h21;
  header[439] = 8'h31;
  header[440] = 8'h06;
  header[441] = 8'h12;
  header[442] = 8'h41;
  header[443] = 8'h51;
  header[444] = 8'h07;
  header[445] = 8'h61;
  header[446] = 8'h71;
  header[447] = 8'h13;
  header[448] = 8'h22;
  header[449] = 8'h32;
  header[450] = 8'h81;
  header[451] = 8'h08;
  header[452] = 8'h14;
  header[453] = 8'h42;
  header[454] = 8'h91;
  header[455] = 8'hA1;
  header[456] = 8'hB1;
  header[457] = 8'hC1;
  header[458] = 8'h09;
  header[459] = 8'h23;
  header[460] = 8'h33;
  header[461] = 8'h52;
  header[462] = 8'hF0;
  header[463] = 8'h15;
  header[464] = 8'h62;
  header[465] = 8'h72;
  header[466] = 8'hD1;
  header[467] = 8'h0A;
  header[468] = 8'h16;
  header[469] = 8'h24;
  header[470] = 8'h34;
  header[471] = 8'hE1;
  header[472] = 8'h25;
  header[473] = 8'hF1;
  header[474] = 8'h17;
  header[475] = 8'h18;
  header[476] = 8'h19;
  header[477] = 8'h1A;
  header[478] = 8'h26;
  header[479] = 8'h27;
  header[480] = 8'h28;
  header[481] = 8'h29;
  header[482] = 8'h2A;
  header[483] = 8'h35;
  header[484] = 8'h36;
  header[485] = 8'h37;
  header[486] = 8'h38;
  header[487] = 8'h39;
  header[488] = 8'h3A;
  header[489] = 8'h43;
  header[490] = 8'h44;
  header[491] = 8'h45;
  header[492] = 8'h46;
  header[493] = 8'h47;
  header[494] = 8'h48;
  header[495] = 8'h49;
  header[496] = 8'h4A;
  header[497] = 8'h53;
  header[498] = 8'h54;
  header[499] = 8'h55;
  header[500] = 8'h56;
  header[501] = 8'h57;
  header[502] = 8'h58;
  header[503] = 8'h59;
  header[504] = 8'h5A;
  header[505] = 8'h63;
  header[506] = 8'h64;
  header[507] = 8'h65;
  header[508] = 8'h66;
  header[509] = 8'h67;
  header[510] = 8'h68;
  header[511] = 8'h69;
  header[512] = 8'h6A;
  header[513] = 8'h73;
  header[514] = 8'h74;
  header[515] = 8'h75;
  header[516] = 8'h76;
  header[517] = 8'h77;
  header[518] = 8'h78;
  header[519] = 8'h79;
  header[520] = 8'h7A;
  header[521] = 8'h82;
  header[522] = 8'h83;
  header[523] = 8'h84;
  header[524] = 8'h85;
  header[525] = 8'h86;
  header[526] = 8'h87;
  header[527] = 8'h88;
  header[528] = 8'h89;
  header[529] = 8'h8A;
  header[530] = 8'h92;
  header[531] = 8'h93;
  header[532] = 8'h94;
  header[533] = 8'h95;
  header[534] = 8'h96;
  header[535] = 8'h97;
  header[536] = 8'h98;
  header[537] = 8'h99;
  header[538] = 8'h9A;
  header[539] = 8'hA2;
  header[540] = 8'hA3;
  header[541] = 8'hA4;
  header[542] = 8'hA5;
  header[543] = 8'hA6;
  header[544] = 8'hA7;
  header[545] = 8'hA8;
  header[546] = 8'hA9;
  header[547] = 8'hAA;
  header[548] = 8'hB2;
  header[549] = 8'hB3;
  header[550] = 8'hB4;
  header[551] = 8'hB5;
  header[552] = 8'hB6;
  header[553] = 8'hB7;
  header[554] = 8'hB8;
  header[555] = 8'hB9;
  header[556] = 8'hBA;
  header[557] = 8'hC2;
  header[558] = 8'hC3;
  header[559] = 8'hC4;
  header[560] = 8'hC5;
  header[561] = 8'hC6;
  header[562] = 8'hC7;
  header[563] = 8'hC8;
  header[564] = 8'hC9;
  header[565] = 8'hCA;
  header[566] = 8'hD2;
  header[567] = 8'hD3;
  header[568] = 8'hD4;
  header[569] = 8'hD5;
  header[570] = 8'hD6;
  header[571] = 8'hD7;
  header[572] = 8'hD8;
  header[573] = 8'hD9;
  header[574] = 8'hDA;
  header[575] = 8'hE2;
  header[576] = 8'hE3;
  header[577] = 8'hE4;
  header[578] = 8'hE5;
  header[579] = 8'hE6;
  header[580] = 8'hE7;
  header[581] = 8'hE8;
  header[582] = 8'hE9;
  header[583] = 8'hEA;
  header[584] = 8'hF2;
  header[585] = 8'hF3;
  header[586] = 8'hF4;
  header[587] = 8'hF5;
  header[588] = 8'hF6;
  header[589] = 8'hF7;
  header[590] = 8'hF8;
  header[591] = 8'hF9;
  header[592] = 8'hFA;
  header[593] = 8'hFF;
  header[594] = 8'hDA;
  header[595] = 8'h00;
  header[596] = 8'h0C;
  header[597] = 8'h03;
  header[598] = 8'h01;
  header[599] = 8'h00;
  header[600] = 8'h02;
  header[601] = 8'h11;
  header[602] = 8'h03;
  header[603] = 8'h11;
  header[604] = 8'h00;
  header[605] = 8'h3F;
  header[606] = 8'h00;
end
